module FP_adder(


);


endmodule

module FP_multiplier(


);

endmodule
